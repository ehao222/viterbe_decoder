`include "params.v"
/*-----------------------------------
// Module: MMU
// File : mmu.v
// Description : Description of MMU Unit in Viterbi Decoder
// Function: used for manage the RAM storing Survivoral Path.
@1.Generate w/r clock
@2 Read Address {ACSPage,ACSSegment};
@3 Read the SurviorBit(8 bit)
@4 Write the stored  SurviorBit(8 bit)
// Simulator : Modelsim 6.5 / Windows 7/10 
-----------------------------------*/
// Revision Number : 1
// Description : Initial Design
/*-----------------------------------*/
module MMU (CLOCK, Clock1, Clock2, Reset, Active, Hold, Init, ACSPage, 
           ACSSegment_minusLSB, Survivors,DataTB, AddressTB,
           RWSelect, ReadClock, WriteClock, RAMEnable, AddressRAM, DataRAM);
// Control
input CLOCK, Clock1, Clock2, Reset, Active, Hold, Init; 
input [`WD_DEPTH-1:0] ACSPage;//the width (6 bit )of theDepth of Tracing back
input [`WD_FSM-2:0] ACSSegment_minusLSB;//5 bit . 256/8=2^5.
// ACS
input [`N_ACS-1:0] Survivors;//4 Survival bits during a clock period.
// TBU
output [`WD_RAM_DATA-1:0] DataTB;//8 bit Survival bits that the Ram Writes
input [`WD_RAM_ADDRESS-`WD_FSM-1:0] AddressTB;//5 bit . 256/8=2^5.
// RAM
output RWSelect, ReadClock, WriteClock, RAMEnable; //RAM W/R control
output [`WD_RAM_ADDRESS-1:0] AddressRAM; //11 bit Address bus
inout [`WD_RAM_DATA-1:0] DataRAM;
//variables
wire [`WD_RAM_DATA-1:0] WrittenSurvivors;//buffer. stores the (4 survival bits*2)=8 bits
reg dummy, SurvRDY;//Period_dummy=(Clock1)*2,Period_SurvRDY=(Clock2)*2,
reg [`WD_RAM_ADDRESS-1:0] AddressRAM; 
reg [`WD_DEPTH-1:0] TBPage;//i.e. Tracking pack depth
wire [`WD_DEPTH-1:0] TBPage_;//TBPage Minus
wire [`WD_DEPTH-1:0] ACSPage;
wire [`WD_TB_ADDRESS-1:0] AddressTB;

initial begin
  dummy<=0;
  SurvRDY<=0;
end
// Read and Write clock
// Dummy variable used because Write Clock only occur every 2 Clocks. 
always @(posedge Clock2 or negedge Reset)
  if (~Reset) dummy <= 0;
  else if (Active) dummy <= ~dummy;
assign WriteClock = (Active && ~dummy) ? Clock1:0;
assign ReadClock = (Active && ~Hold) ? ~Clock1:0; 
// For Survivor Buffer,
// -- The buffer used because Data Bus Width is 8, while
// ACS output is only 4 bits at one time
always @(posedge Clock1 or negedge Reset)
  if (~Reset) SurvRDY <= 1; 
  else if (Active) SurvRDY <= ~SurvRDY;
ACSSURVIVORBUFFER buff (Reset, Clock1, Active, SurvRDY, Survivors,
             WrittenSurvivors);
// --
// For Traceback Ops
// every negedge Clock2 : - TBPage is decreased by 1, OR
// - When Init is Active, TBPage equal ACSPage - 1 
always @(negedge Clock2 or negedge Reset)begin
  if (~Reset) begin 
  TBPage <= 0;
  end
  else if (Init) TBPage <= ACSPage-1;
  else TBPage <= TBPage_;
end

assign TBPage_ = TBPage - 1;
assign RAMEnable = 0;
assign RWSelect = (Clock2) ? 1:0;//RWSelect=Clock2
assign DataRAM = (~Clock2) ? WrittenSurvivors:'bz; //(0:ACS->RAM)
assign DataTB = (Clock2) ? DataRAM:'bz;//(1:RAM->TBU)
// every time Clock2 changes, the Address and Enable for each RAM has to
// be set so it will be ready when Read/Write Clock occur on the edges of // Clock1.
always @(posedge CLOCK or negedge Reset)begin
  if (~Reset) AddressRAM <= 0;
  else if (Active) begin
      if (Clock2 == 0) // this is when read happened begin
      AddressRAM <= {ACSPage, ACSSegment_minusLSB}; 
  end
  else 
    AddressRAM <= {TBPage [`WD_DEPTH-1:0],AddressTB};  
  end
//--
endmodule

/*-----------------------
//Module:ACSSURVIVORBUFFER
// File : mmu.v
// Description :
-----------------------*/
/*-----------------------------------*/
module ACSSURVIVORBUFFER (Reset, Clock1, Active, SurvRDY, Survivors,
WrittenSurvivors);
/*-----------------------------------------
//Clock1
//SurvRDY:Div2_CLOCK1
//Survivors: 4-bits survival bits generated by ACS
//WrittenSurvivors:8-bits survival bits 
// To accomodate the use of 8 bit wide RAM DATA BUS, the Survivor
// (which is only 4 on every clock) must be buffered first.

            | Surviors        |
            |   /|\           | 
Survivors ->| WrittenSurviors_|<=>WrittenSurviors
            |                 |
-----------------------------------------*/
input Reset, Clock1, Active, SurvRDY;
input [`N_ACS-1:0] Survivors;
output [`WD_RAM_DATA-1:0] WrittenSurvivors;
wire [`WD_RAM_DATA-1:0] WrittenSurvivors;
reg [`N_ACS-1:0] WrittenSurvivors_;//low 4 bits
always @(posedge Clock1 or negedge Reset) begin
  if (~Reset) WrittenSurvivors_ = 0; 
  else if (Active)
    WrittenSurvivors_ = Survivors; 
end
assign WrittenSurvivors = (SurvRDY) ? {Survivors, WrittenSurvivors_}:8'bz; 
endmodule