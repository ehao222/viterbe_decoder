`include "params.v"
/*-----------------------------------*/
// Module: VITERBIDECODER
// File : decoder.v
// Description : Top Level Module of Viterbi Decoder 
// Simulator : Modelsim 6.5 / Windows 7/10 
/*-----------------------------------*/
// Revision Number : 1
// Description : Initial Design 
/*-----------------------------------*/
//module VITERBIDECODER (Reset, CLOCK, Active, Code, DecodeOut); 
module VITERBIDECODER (Reset, CLOCK, Active, Code, DecodeOut);
//复位，时钟，激活标志位，解码输出
input Reset, CLOCK, Active; 
input [`WD_CODE-1:0] Code;//解码输入 ，位宽为2
output DecodeOut;
wire [`WD_DIST*2*`N_ACS-1:0] Distance; // BMG Output 计算位宽：16=分支度量宽度*分支数*4个状态
wire [`WD_FSM-1:0] ACSSegment; //处理后的状态段，4个ACS，共256个状态，需要迭代64次迭代
wire [`WD_DEPTH-1:0] ACSPage; //control输出
wire CompareStart, Hold, Init;//CompareStart标志加比选模块是否进行比较操作，对于第一个(K-1)进程，在每个节点上只有一个输入
wire [`N_ACS-1:0] Survivors;//acs输出
wire [`WD_STATE-1:0] LowestState;//幸存信息比特*4
wire TB_EN;//最小路径度量状态
wire RAMEnable;
wire ReadClock, WriteClock, RWSelect;
wire [`WD_RAM_ADDRESS-1:0] AddressRAM;// RAM AddressBus, // generated by TBU and ACSURAM 地址总线
wire [`WD_RAM_DATA-1:0] DataRAM; // RAM Databus ，RAM 数据总线
wire [`WD_RAM_DATA-1:0] DataTB;
wire [`WD_RAM_ADDRESS-`WD_FSM-1:0] AddressTB; 
wire Clock1, Clock2;
// for metric memory connection 度量内存连接 
wire [`WD_METR*2*`N_ACS-1:0] MMPathMetric; //内存读取的路径度量(old)64bit
wire [`WD_METR*`N_ACS-1:0] MMMetric;//路径度量，Metric-->MMMetric
wire [`WD_FSM-2:0] MMReadAddress;//读地址：5bit位宽
wire [`WD_FSM-1:0] MMWriteAddress;//内存接口写地址6bit
wire MMBlockSelect;//存储块选：1bit
// instantiation of Viterbi Decoder Modules 维特比译码器模块的实例化 
CONTROL ctl (Reset, CLOCK, Clock1, Clock2, ACSPage, ACSSegment,Active, CompareStart, Hold, Init, TB_EN);
BMG bmg (Reset, Clock2, ACSSegment, Code, Distance);
ACSUNIT acs (Reset, Clock1, Clock2, Active, Init, Hold, CompareStart, ACSSegment,
     Distance, Survivors, LowestState,MMReadAddress, MMWriteAddress, MMBlockSelect, 
     MMMetric, MMPathMetric);

MMU mmu (CLOCK, Clock1, Clock2, Reset, Active, Hold, Init, ACSPage, 
     ACSSegment [`WD_FSM-1:1], Survivors,DataTB, AddressTB,RWSelect,
      ReadClock, WriteClock, RAMEnable, AddressRAM, DataRAM);

TBU tbu (Reset, Clock1, Clock2, TB_EN, Init, Hold, LowestState, 
        DecodeOut, DataTB, AddressTB);

METRICMEMORY mm (Reset, Clock1, Active, MMReadAddress, MMWriteAddress, 
      MMBlockSelect, MMMetric, MMPathMetric);

RAM ram (RAMEnable, AddressRAM, DataRAM, RWSelect, ReadClock, WriteClock); 
endmodule